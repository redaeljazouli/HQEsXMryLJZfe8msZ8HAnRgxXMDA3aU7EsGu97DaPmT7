compteur60_inst : compteur60 PORT MAP (
		aclr	 => aclr_sig,
		aset	 => aset_sig,
		clock	 => clock_sig,
		cnt_en	 => cnt_en_sig,
		updown	 => updown_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
